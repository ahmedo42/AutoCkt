cs_amp test
.include "/home/ksettaluri6/AutoCkt/eval_engines/ngspice/ngspice_inputs/spice_models/45nm_bulk.txt"

.param  vbias=0.8
.param  rload=500
.param  cload=100f
.param  mul=12
.param  L=0.18u E=0.54u W=0.8u  as="W*E"    ad="W*E"    ps="2*(E+W)"    pd="2*(E+W)"

M1  vd  vg  0   0   NMOS  w=W    l=L  as=as   ad=ad   ps=ps   PD=pd  m=mul

Rl  VDD vd  rload
Cl  vd  0   cload

Vdd VDD 0   1.8
vin vg  0   dc=vbias    ac=1

.ac dec 20  1Meg  100G

.control
run
set wr_vecnames
option numdgt=7
wrdata ac.csv vm(vd)
op
wrdata dc.csv i(Vdd)
.endc

.end